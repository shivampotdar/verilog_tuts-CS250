// 4 bit RCA

module TB_RCA_4b();

    // internal vars
    reg [3:0] A, B;   /* A and B are 4 elements */
    /* input [3:0] A[3:0] means every element of A is 4b array*/
    reg carry_in;
    wire [3:0] Sum;
    wire carry_out;

    // instantiate

    RCA_4b rca_4b_dut(Sum, carry_out, A, B, carry_in);

    initial
    begin
        
        $monitor($time,".A : %d B : %d carry_in : %b Sum : %d carry_out : %b",A,B,carry_in,Sum,carry_out);
        $dumpsfile("TB_RCA_4b.vcd");
        $dumpvars(0,TB_RCA_4b);
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 0; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 0; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 0; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 0; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 0; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 0; B[1]= 1; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 0; B[0]= 1; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 0; carry_in= 1;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 0;
#5  A[3]= 1; A[2]= 1; A[1]= 1; A[0]= 1; B[3]= 1; B[2]= 1; B[1]= 1; B[0]= 1; carry_in= 1;


end

endmodule
